// Code your design here
`include"ALU.sv"
`include"Ctrl.sv"
`include"DMem.sv"
`include"InstROM.sv"
`include"JLUT.sv"
`include"ProgCtr.sv"
`include"RegFile.sv"
`include"Top.sv"